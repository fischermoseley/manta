../../../common/divider.sv