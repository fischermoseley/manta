/*
This playback module was generated with Manta /* VERSION */ on /* TIMESTAMP */ by /* USER */

If this breaks or if you've got dank formal verification memes, contact fischerm [at] mit.edu

Provided under a GNU GPLv3 license. Go wild.

Here's an example instantiation of the Manta module you configured, feel free to copy-paste
this into your source!

manta manta_inst (
    .clk(clk),

    /* EX_INST_PORTS */);

*/

module manta(
    input wire clk,

    /* TOP_LEVEL_PORTS */);


    /* INTERFACE_RX */

    /* CORE_CHAIN */

    /* INTERFACE_TX */

endmodule

/* ---- Module Definitions ----  */

/* MODULE_DEFS */