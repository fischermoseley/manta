`default_nettype none
`timescale 1ns / 1ps

module top_level (
	input wire clk,

    output logic [15:0] led,
    output logic ca, cb, cc, cd, ce, cf, cg,
    output logic [7:0] an,

    output logic led16_r,
    output logic led17_r,

    output reg eth_refclk,
    output reg eth_rstn,

    input wire eth_crsdv,
    input wire [1:0] eth_rxd,

    output reg eth_txen,
    output reg [1:0] eth_txd);

    assign eth_rstn = 1;

    logic clk_50mhz;
    assign eth_refclk = clk_50mhz;
    divider d (.clk(clk), .ethclk(clk_50mhz));

    assign led = manta_inst.brx_my_lut_ram_addr;
    assign led16_r = manta_inst.brx_my_lut_ram_rw;
    assign led17_r = manta_inst.brx_my_lut_ram_valid;

    ssd ssd (
        .clk(clk_50mhz),
        .val( {manta_inst.my_lut_ram_btx_rdata, manta_inst.brx_my_lut_ram_wdata} ),
        .cat({cg,cf,ce,cd,cc,cb,ca}),
        .an(an));

    manta manta_inst (
        .clk(clk_50mhz),

        .crsdv(eth_crsdv),
        .rxd(eth_rxd),
        .txen(eth_txen),
        .txd(eth_txd));


endmodule

`default_nettype wire